class transaction;
  
  bit [31:0] concatenated;
  
  bit [7:0] button_counter;
  
endclass