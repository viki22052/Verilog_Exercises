class transaction;
  
  bit btn;
  
  bit [7:0] button_counter;
  
endclass