
module andFunct(a, b, out);
input a, b;
output out;
wire out = a & b;

endmodule

