interface bct_tb(input logic clk, rst);
  
  logic [31:0] concatenated;
  logic [7:0] button_counter;
  
  
  
  
endinterface 