interface bct_tb(input logic clk, rst);
  
  logic btn;
  logic [7:0] button_counter;
  
  
  
  
endinterface 